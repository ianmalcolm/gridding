`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:26:10 07/06/2016 
// Design Name: 
// Module Name:    GRIDDING 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module GRIDDING(
    input [31:0] sampleDataR,
    input [31:0] sampleDataI,
    input [31:0] sampleIu,
    input [31:0] sampleIv,
    input [31:0] sampleOffset,
    input clk,
    input rst,
    input [31:0] addr,
    output [31:0] data
    );


endmodule
